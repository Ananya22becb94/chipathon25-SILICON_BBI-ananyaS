magic
tech gf180mcuD
timestamp 1678205252
<< nwell >>
rect 0 102 76 166
<< nmos >>
rect 16 21 22 38
rect 33 21 39 38
rect 50 21 56 38
<< pmos >>
rect 19 111 25 145
rect 30 111 36 145
rect 50 111 56 145
<< ndiff >>
rect 6 36 16 38
rect 6 23 8 36
rect 13 23 16 36
rect 6 21 16 23
rect 22 36 33 38
rect 22 23 25 36
rect 30 23 33 36
rect 22 21 33 23
rect 39 36 50 38
rect 39 23 42 36
rect 47 23 50 36
rect 39 21 50 23
rect 56 36 66 38
rect 56 23 59 36
rect 64 23 66 36
rect 56 21 66 23
<< pdiff >>
rect 9 143 19 145
rect 9 113 11 143
rect 16 113 19 143
rect 9 111 19 113
rect 25 111 30 145
rect 36 143 50 145
rect 36 113 39 143
rect 47 113 50 143
rect 36 111 50 113
rect 56 143 66 145
rect 56 113 59 143
rect 64 113 66 143
rect 56 111 66 113
<< ndiffc >>
rect 8 23 13 36
rect 25 23 30 36
rect 42 23 47 36
rect 59 23 64 36
<< pdiffc >>
rect 11 113 16 143
rect 39 113 47 143
rect 59 113 64 143
<< psubdiff >>
rect 6 12 21 14
rect 6 7 11 12
rect 16 7 21 12
rect 6 5 21 7
rect 30 12 45 14
rect 30 7 35 12
rect 40 7 45 12
rect 30 5 45 7
rect 54 12 69 14
rect 54 7 59 12
rect 64 7 69 12
rect 54 5 69 7
<< nsubdiff >>
rect 6 159 21 161
rect 6 154 11 159
rect 16 154 21 159
rect 6 152 21 154
rect 30 159 45 161
rect 30 154 35 159
rect 40 154 45 159
rect 30 152 45 154
rect 54 159 69 161
rect 54 154 59 159
rect 64 154 69 159
rect 54 152 69 154
<< psubdiffcont >>
rect 11 7 16 12
rect 35 7 40 12
rect 59 7 64 12
<< nsubdiffcont >>
rect 11 154 16 159
rect 35 154 40 159
rect 59 154 64 159
<< polysilicon >>
rect 19 145 25 150
rect 30 145 36 150
rect 50 145 56 150
rect 19 107 25 111
rect 16 102 25 107
rect 30 108 36 111
rect 30 102 39 108
rect 16 80 22 102
rect 16 78 28 80
rect 16 72 20 78
rect 26 72 28 78
rect 16 70 28 72
rect 16 38 22 70
rect 33 67 39 102
rect 50 93 56 111
rect 44 91 56 93
rect 44 85 46 91
rect 52 85 56 91
rect 44 83 56 85
rect 33 65 43 67
rect 33 59 35 65
rect 41 59 43 65
rect 33 57 43 59
rect 33 38 39 57
rect 50 38 56 83
rect 16 16 22 21
rect 33 16 39 21
rect 50 16 56 21
<< polycontact >>
rect 20 72 26 78
rect 46 85 52 91
rect 35 59 41 65
<< metal1 >>
rect 0 159 76 166
rect 0 154 11 159
rect 16 154 35 159
rect 40 154 59 159
rect 64 154 76 159
rect 0 152 76 154
rect 11 143 16 145
rect 11 112 16 113
rect 8 107 16 112
rect 39 143 47 152
rect 39 111 47 113
rect 59 143 64 145
rect 8 91 13 107
rect 59 104 64 113
rect 59 98 61 104
rect 67 98 69 104
rect 8 85 46 91
rect 52 85 54 91
rect 8 51 13 85
rect 18 72 20 78
rect 26 72 28 78
rect 33 59 35 65
rect 41 59 43 65
rect 8 46 30 51
rect 8 36 13 38
rect 8 14 13 23
rect 25 36 30 46
rect 25 21 30 23
rect 42 36 47 38
rect 42 14 47 23
rect 59 36 64 98
rect 59 21 64 23
rect 0 12 76 14
rect 0 7 11 12
rect 16 7 35 12
rect 40 7 59 12
rect 64 7 76 12
rect 0 0 76 7
<< via1 >>
rect 61 98 67 104
rect 46 85 52 91
rect 20 72 26 78
rect 35 59 41 65
<< metal2 >>
rect 59 104 69 105
rect 59 98 61 104
rect 67 98 69 104
rect 59 97 69 98
rect 44 91 54 92
rect 44 85 46 91
rect 52 85 54 91
rect 44 84 54 85
rect 18 78 28 79
rect 18 72 20 78
rect 26 72 28 78
rect 18 71 28 72
rect 33 65 43 66
rect 33 59 35 65
rect 41 59 43 65
rect 33 58 43 59
<< labels >>
rlabel metal2 23 75 23 75 1 A
port 1 n
rlabel metal2 38 62 38 62 1 B
port 2 n
rlabel metal2 64 101 64 101 1 Y
port 3 n
rlabel nsubdiffcont 13 156 13 156 1 VDD
port 4 n
rlabel psubdiffcont 13 9 13 9 1 VSS
port 5 n
<< end >>
